`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/09/30 12:20:06
// Design Name: 
// Module Name: top_7seg_demo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module top_7seg_demo(CLK100MHZ,reset,CA,CB,CC,CD,CE,CF,CG, AN );
input CLK100MHZ, reset;
output CA, CB,CC,CD,CE,CF,CG;
output [7:0] AN;   
wire en;
wire [3:0] D0,D1,D2,D3,D4,D5,D6,D7;

seven_segement_8_drv u0 (.clk(CLK100MHZ), .reset(!reset),.D0(D0), .D1(D1), .D2(D2), .D3(D3),
                        .D4(D4), .D5(D5), .D6(D6), .D7(D7), .a(CA), .b(CB), .c(CC), .d(CD), 
                        .e(CE), .f(CF), .g(CG),.AN(AN));
                        
bcd_cnt cnt(.Q(D0), .TC(), .inc(en), .rstn(!reset), .clk(CLK100MHZ));
cnt_100M div(.clk(CLK100MHZ), .rstn(!reset), .eo_100M(en), .eo_10k(), .eo_1k()); 

assign D1 = D0+1;   
assign D2 = D0+2;  
assign D3 = D0+3; 
assign D4 = D0+4; 
assign D5 = D0+5; 
assign D6 = D0+6; 
assign D7 = D0+7;
 
endmodule
